

module decoder
    #(
		parameter A_SIZE = 3,	// ALU function width
		parameter O_SIZE = 6	// OpCode width
    )
    (
		// Outputs
		output cpuConfig::aluFunc_t aluFunc,
		output logic aluImmediate,
		output logic immSwitches,
		output logic pcInc,
		output logic writeReg,

		input cpuConfig::opCode_t opCode,
		input wire demoSwitch
	);
	

	import cpuConfig::*;


	always_comb begin
		// Set default values
		aluFunc = ALU_A;
		aluImmediate = 1'b0;
		immSwitches = 1'b0;
		pcInc = 1'b1;
		writeReg = 1'b1;

		// Decode opCode
		case (opCode)
			LDI: begin
				aluFunc = ALU_B;
				aluImmediate = 1'b1;
			end
			LDS: begin
				pcInc = demoSwitch;

				aluFunc = ALU_B;
				aluImmediate = 1'b1;
				immSwitches = 1'b1;
			end
			ADD: begin
				aluFunc = ALU_ADD;
			end
			ADDI: begin
				aluFunc = ALU_ADD;
				aluImmediate = 1'b1;
			end
			MUL: begin
				aluFunc = ALU_MUL;
			end
			MULI: begin
				aluFunc = ALU_MUL;
				aluImmediate = 1'b1;
			end
			WAIT0: begin
				pcInc = ~demoSwitch;
			end
			WAIT1: begin
				pcInc = demoSwitch;
			end
		endcase
	end


endmodule
