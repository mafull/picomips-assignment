'define F_SIZE 2

'define 