module registers
    #(

    )
    (

    );


endmodule
